`define BASE 5
`define LOGBASE 3
`define DIGITWIDTH 3
`define SEQWIDTH 7

// `define DIGITWIDTH 4
// `define SEQWIDTH 9
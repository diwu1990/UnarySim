`define GCWD 8
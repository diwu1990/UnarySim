`define BASE 2
`define LOGBASE 1
`define DIGITWIDTH 8
`define SEQWIDTH 8
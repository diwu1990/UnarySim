`define BASE 3
`define LOGBASE 2
`define DIGITWIDTH 5
`define SEQWIDTH 8

// `define DIGITWIDTH 3
// `define SEQWIDTH 6
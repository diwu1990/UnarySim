`include "SobolSeq2Def.sv"
module SobolSeq2 (
    input logic clk,    // Clock
    input logic rst,  // Asynchronous reset active low
    input logic in,
    input logic out
);

endmodule
`define GWIDTH 4
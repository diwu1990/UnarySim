`ifndef MAC_BW
    `define MAC_BW 8
`endif

`ifndef MAC_CNT
    `define MAC_CNT 16
`endif

`ifndef ROW_CNT
    `define ROW_CNT 16
`endif

`ifndef COL_CNT
    `define COL_CNT 16
`endif

`ifndef ADDR_BW
    `define ADDR_BW 4
`endif
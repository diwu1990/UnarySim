`define INWIDTH 8
`define LOGINWIDTH 3
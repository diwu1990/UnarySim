`define INWD 8
`define LOGINWD 3
